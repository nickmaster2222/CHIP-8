import types::*;
package imports;

typedef struct {
	u8 opcode,
	u5 r1,
	u5 r2,
	u8 val1,
	u8 val2,
	u16 I
} chip8_instruction;



endpackage